`ifndef PKT_GEN_SV
`define PKT_GEN_SV


`endif